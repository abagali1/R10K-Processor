/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  branch_fu_test.sv                                   //
//                                                                     //
//  Description :  Testbench module for the branch FU                  //
//                                                                     //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`include "sys_defs.svh"
`include "ISA.svh"