`include "sys_defs.svh"

